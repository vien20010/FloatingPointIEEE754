`timescale 1ns / 1ps
`include "add_sub.sv"

module add_sub_tb;
	logic 	[31:0]	A,B;
	logic	[31:0]	result;
	logic 			underflag,overflag;

	
	logic				add_or_sub;


	add_sub uut(.A(A),
				.B(B),
				.checkequation(add_or_sub),
				.overflow(overflag),
				.underflow(underflag),
				.result(result));

	initial
		begin
				add_or_sub = 1;
				
    A = 32'b01000000101000000000000000000000;
    B = 32'b01000000111000000000000000000000;
    
    #10;
    A = 32'b01000000101000000000000000000000;
    B = 32'b01000000111000000000000000000000;

    #10;
    A = 32'b11000001011110011001100110011010; //-15.6
    B = 32'b01000000011011001100110011001101; // 3.7

    #10;
    A = 32'b11000001011110011001100110011010; //-15.6
    B = 32'b01000000011011001100110011001101; // 3.7

    #10;
    A = 32'b11000001011110011001100110011010; // 15.6
    B = 32'b11000000011011001100110011001101; // 3.7

    #10;
    A = 32'b11000000111100001111010111000011; // -7.53
    B = 32'b01000011010101111001010001111011; // 215.58

    #10;
    A = 32'b11000000111100001111010111000011; // -7.53
    B = 32'b01000011010101111001010001111011; // 215.58

    #10;
    A = 32'b00111100101101011101110011000110; //0.0222 
    B = 32'b00111111011010001111010111000011; //0.91

    #10;
    B = 32'b00111100101101011101110011000110; //0.0222 
    A = 32'b00111111011010001111010111000011; //0.91

    #10;
    A = 32'b01111111100000000000000000000000; // Inf
    B = 32'b01000000011011001100110011001101; // 3.7

    #10;
    A = 32'b01111111100000000000000000000000; // Inf
    B = 32'b01000000011011001100110011001101; // 3.7

    #10;
    A = 32'b01111111100000000000000000000000; // Inf
    B = 32'b01111111100000000000000000000000; // Inf

    #10;
    A = 32'b11111111100000000000000000000000; // -Inf
    B = 32'b11111111100000000000000000000000; // -Inf

    #10;
    A = 32'b01111111100000000000000000000000; // +Inf
    B = 32'b11111111100000000000000000000000; // -Inf

    #10;
    A = 32'b11111111100000000000000000000000; // -Inf
    B = 32'b01111111100000000000000000000000; // +Inf

    #10;
    A = 32'b11111111100000000000000000000000; // -Inf
    B = 32'b01111111100000000000000000000000; // +Inf


    #10;
    A = 32'b01111111100000000000000000000000; // Inf
    B = 32'b01111111100000000000000000000000; // Inf

    #10;
    A = 32'b11111111100000000000000000000000; // -Inf
    B = 32'b11111111100000000000000000000000; // -Inf

    #10;
    A = 32'b01111111100000000000000000000000; // +Inf
    B = 32'b11111111100000000000000000000000; // -Inf

    #10;
    A = 32'b11111111100000000000000000000000; // -Inf
    B = 32'b01111111100000000000000000000000; // +Inf

    #10;
    A = 32'b11111111100000000000000000000000; // -Inf
    B = 32'b01111111100000000000000000000000; // +Inf

    #10;
    A = 32'b01111111100000000000000000000000; // Inf
    B = 32'b11111111100000000000000000000001; // NaN

    #10;
    A = 32'b10111111011010100000011010001111; //-0.9141625863
    B = 32'b00111011000100011010001010110100; //0.00222222222

    #10;
    A = 32'b00000000000000000000000000000000; // 0
    B = 32'b01000000011011001100110011001101; // 3.7

    #10;
    A = 32'b01000000011011001100110011001101; // 3.7
    B = 32'b01000000011011001100110011001101; // 3.7

    #10;
    A = 32'b00000000000000000000000000000000; // 3.7
    B = 32'b01000000011011001100110011001101; // 3.7

    #10;
    A = 32'b01111111100000000000000000000000; // Inf
    B = 32'b01000000011011001100110011001101; // 3.7

    #10;
    A = 32'b01111111100000000000000000000000; // Inf
    B = 32'b11111111100000000000000000000001; // NaN

    #10;

    // Long Add // Failed case
    A = 32'b00111111100000100000100000010111; // 
    B = 32'b00110101001011101011100111101101; // 

    #10;
    A = 32'b00111111011111111110011011100111; // 
    B = 32'b10101101001001001110011011110010; // 

    #10;
    A = 32'b00111111011111111110100010001101; // 
    B = 32'b10101101000001100111001000101101; // 

    #10;
    A = 32'b00111111011111111101011011010001; // 
    B = 32'b10101110001101100010010001010001; // 

    #10;
			
			$finish;
		end

endmodule
