`timescale 1ns / 1ps
`include "mult.sv"
`include "mult24_booth.sv"
`include "adder.sv"
`include "sub.sv"
`include "find1.sv"
`include "complement2.sv"
`include "shiftleft24.sv"
`include "shiftleft48.sv"
`include "shift_right.sv"
`include "export_result.sv"
`include "checkspecial.sv"


module multiplier_tb;
logic [31:0]A,B;
   logic [31:0]result;
    logic underflow,overflow;

    


    mult uut(.A(A),
                .B(B),
                .overflow(overflow),
                .underflow(underflow),
                .result(result));

initial begin
	A = 32'b01000000000000000000000000000000;

	B = 32'b00111111100000000000000000000000;
	#50;

	A = 32'b01000000000000000000000000000000;

	B = 32'b01000000000000000000000000000000;
	#50;
	
	A = 32'b01000000101010000000000000000000;

	B = 32'b01000000000000000000000000000000;
	#50;
	A = 32'b10111111100000000000000000000000; //-1

	B = 32'b01000000000000000000000000000000;
	#50;
	A = 32'b01000000001000000000000000000000; //2.5

	B = 32'b01000000011000000000000000000000; //3.5
	#50;
	A = 32'b01000100111111000111001100110011; //2019.6
	
	B = 32'b11000000011000000000000000000000; //-3.5
	#50;

	A = 32'b01000100111111000111001100110011; //2019.6
	
	B = 32'b11111111100000000000000000000001;// NaN

	#50;
	A = 32'b0_00000000_00000000000000000000000; // 0
	
	B = 32'b0_00000000_00000000000000000000000; // 0

	#50;
	A = 32'b1_11111111_00000000000000000000000;// -INF
	
	B = 32'b0_11111111_00000000000000000000000;// +INF

	#50;
	A = 32'b0_11111111_00000000000000000000000;// +INF
	
	B = 32'b0_00000000_00000000000000000000000;// 0

	#50;
	A = 32'b1_11111111_00000000000000000000000;// -INF
	
	B = 32'b1_11111111_00000000000000000000000;// -INF

	#50;
	A = 32'b0_11111111_00000000000000000000000;// +INF
	
	B = 32'b1_11111111_00000000000000000000000;// -INF

	A = 32'b00111101100000100000100000010111; // 
	B = 32'b00110101001011101011100111101101; // 
	#50;
	A = 32'b00111011011111111110011011100111; // 
	B = 32'b10101101001001001110011011110010; // 
	#50;
	A = 32'b00110111011111111110100010001101; // 
	B = 32'b10101101000001100111001000101101; // 
	#50;
	A = 32'b00101111011111111101011011010001; // 
	B = 32'b10101110001101100010010001010001; // 
	#50;
	$finish;

end

endmodule