

module TAYLOR_EXP_tb();

logic [31:0] in;
logic [31:0] out;


TAYLOR_EXP TAYLOR_EXP_0 (.in(in),.out(out));

initial begin
	
	
	#10
	in = 32'b00111010100000110001001001101111; // 0.001
	#10
	in = 32'b00111100001000111101011100001010; // 0.01
	#10
	in = 32'b00111101110011001100110011001101; // 0.1
	#10
    in = 32'b01000001001000000000000000000000; // 10
    #10
    in = 32'b01000000000000000000000000000000; // 2
    #10
    in = 32'b00111111110000111101011100001010; // 1.53
	#10
    in = 32'b00111111000001101010011111110000; // 0.526
    #10
    in = 32'b10111111000001101010011111110000; // -0.526
    #10
    in = 32'b10111111110000111101011100001010; // -1.53
	
end


endmodule 